package myPackage;
    module a();
    endmodule

endpackage